// Copyright 2022 Politecnico di Torino.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 2.0 (the "License"); you may not use this file except in
// compliance with the License. You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-2.0. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// File: fpu_if.sv
// Author: Michele Caon
// Date: 31/05/2022

/*
 * File: fpu_if.sv
 * ----------------------------------------
 * Interface with the fpu wrapper in 'fpu_wrap.sv'.
 */

import fpnew_pkg::*;
import cf_math_pkg::*;

interface fpu_if #();

    /* INTERFACE SIGNALS */
    logic                               clk,
    logic                               rst,
    logic [NUM_OPERANDS-1:0][WIDTH-1:0] operands,
    fpnew_pkg::roundmode_e              rnd_mode,
    fpnew_pkg::operation_e              op,
    logic                               op_mod,
    fpnew_pkg::fp_format_e              src_fmt,
    fpnew_pkg::fp_format_e              dst_fmt,
    fpnew_pkg::int_format_e             int_fmt,
    logic                               vectorial_op,
    TagType                             tag,
    logic                               in_valid,
    logic                               in_ready,
    logic                               flush,
    logic [WIDTH-1:0]                   result,
    fpnew_pkg::status_t                 status,
    TagType                             tag,
    logic                               out_valid,
    logic                               out_ready,
    logic                               busy

    /* INTERFACE SIGNALS MODE MAPPING */

    /* Interface port at ALU side (DUT) */
    modport fpu_port (
        input logic                               clk,
        input logic                               rst,
        input logic [NUM_OPERANDS-1:0][WIDTH-1:0] operands,
        input fpnew_pkg::roundmode_e              rnd_mode,
        input fpnew_pkg::operation_e              op,
        input logic                               op_mod,
        input fpnew_pkg::fp_format_e              src_fmt,
        input fpnew_pkg::fp_format_e              dst_fmt,
        input fpnew_pkg::int_format_e             int_fmt,
        input logic                               vectorial_op,
        input TagType                             tag,
        input logic                               in_valid,
        output logic                               in_ready,
        input logic                               flush,
        output logic [WIDTH-1:0]                  result,
        output fpnew_pkg::status_t                status,
        output TagType                            tag,
        output logic                              out_valid,
        input  logic                              out_ready,
        output logic                              busy   
    );

    /* Interface port at driver side (unused since the driver is a class) */
    modport driver_port (
        output logic                               clk,
        output logic                               rst,
        output logic [NUM_OPERANDS-1:0][WIDTH-1:0] operands,
        output fpnew_pkg::roundmode_e              rnd_mode,
        output fpnew_pkg::operation_e              op,
        output logic                               op_mod,
        output fpnew_pkg::fp_format_e              src_fmt,
        output fpnew_pkg::fp_format_e              dst_fmt,
        output fpnew_pkg::int_format_e             int_fmt,
        output logic                               vectorial_op,
        output TagType                             tag,
        output logic                               in_valid,
        input logic                                in_ready_
        output logic                               flush,
        input logic [WIDTH-1:0]                    result,
        input fpnew_pkg::status_t                  status,
        input TagType                              tag,
        input logic                                out_valid,
        output logic                               out_ready,
        input logic                                busy  
    );

    /*
     * NOTE: an interface can be used to abstract the communication
     * with a module and to implement self-checking functions. In 
     * this case, we use it to generate the clock for the sequential
     * ALU and to check that the result is consistent with the input.
     */

    /******************************************************************************/
    /* CLOCK GENERATION */

    // Initialize clock and reset
    initial begin: init
        clk_i    = 1'b1;
        rst_ni   = 1'b1;
    end

    // Generate clock
    always #5ns begin: clk_gen
        clk_i= ~clk_i
    end

    // Reset the DUT
    task rst_dut();
        @(negedge clk_i;
        rst_ni   = 1'b0;
        @(negedge clk_i;
        rst_ni   = 1'b1;
    endtask // rst_dut

    // ----------
    // ASSERTIONS
    // ----------
    `ifndef SYNTHESIS
    `include "fpu_if_sva.svh"
    `endif /* SYNTHESIS */

endinterface // fpu_if